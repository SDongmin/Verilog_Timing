module led_dir(
	input clk, clk_1k, reset,
	output reg [15:0] led
);

reg [3:0] count;
reg [9:0] c;



end



endmodule
